`ifndef COMMON_DEFS_SVH
`define COMMON_DEFS_SVH

`define INT_BITS    8
`define FRAC_BITS   24
`define WORD_WIDTH   (`INT_BITS+`FRAC_BITS)

`define SCREEN_WIDTH    640
`define SCREEN_HEIGHT   480

`define COLOR_WIDTH     24


`endif // COMMON_DEFS_SVH
